LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE compiled IS
    TYPE binary IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR (15 DOWNTO 0);
END PACKAGE;