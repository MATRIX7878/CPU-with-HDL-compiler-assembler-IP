LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY work;
USE WORK.compiled.ALL;
USE WORK.translator.ALL;

ENTITY CPU_TB IS
END ENTITY;

ARCHITECTURE behavior OF CPU_TB IS

SIGNAL clk : STD_LOGIC := '1';
SIGNAL assembled : STD_LOGIC := '0';
SIGNAL raw : STD_LOGIC_VECTOR (2047 DOWNTO 0) := (OTHERS => '0');
SIGNAL CMD : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
SIGNAL ARG : STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
SIGNAL machine : binary := (OTHERS => (OTHERS => '0'));

BEGIN
	clk <= NOT clk after 18.5 ns;
	raw(2047 DOWNTO 1232) <= x"434C522041430A53544120420A4A4D505A2031300A0A2E6F72672031300A41444420420A41444420310A53544120420A535441204C45440A505345203235300A505345203235300A505345203235300A505345203235300A434C522041430A4A4D505A203130";

	PARSE_int : entity work.parser
		PORT MAP(clk => clk, raw => raw, CMD => CMD, ARG => ARG);
	ASSEMBLER_int : entity work.assembler
		PORT MAP(clk => clk, instruction => CMD, input => ARG, assembled => assembled, machine => machine);
	TOPLEVEL_inst : entity work.toplevel
   		PORT MAP(clk => clk);
END ARCHITECTURE;