PACKAGE flashStates IS
    TYPE state IS (INIT, LOADCMD, LOADADDR, LOADDATA, SEND, READ, DONE);
END PACKAGE;